library ieee;
    use ieee.numeric_std.all;
    use ieee.std_logic_1164.all;

entity DTM_Bscane2 is
    port (
        i_clk : in std_logic
    );
end entity DTM_Bscane2;

architecture rtl of DTM_Bscane2 is
    
begin
    
    
    
end architecture rtl;