library ieee;
    use ieee.numeric_std.all;
    use ieee.std_logic_1164.all;

entity DebugModule is
    port (
        i_clk : in std_logic
    );
end entity DebugModule;

architecture rtl of DebugModule is
    
begin
    
    
    
end architecture rtl;